magic
tech scmos
timestamp 1725621116
<< nwell >>
rect -2 -9 23 12
rect 36 -9 61 12
<< ntransistor >>
rect 9 -21 11 -17
rect 47 -21 49 -17
<< ptransistor >>
rect 9 -2 11 6
rect 47 -2 49 6
<< ndiffusion >>
rect 8 -21 9 -17
rect 11 -21 12 -17
rect 46 -21 47 -17
rect 49 -21 50 -17
<< pdiffusion >>
rect 8 -2 9 6
rect 11 -2 12 6
rect 46 -2 47 6
rect 49 -2 50 6
<< ndcontact >>
rect 4 -21 8 -17
rect 12 -21 16 -17
rect 42 -21 46 -17
rect 50 -21 54 -17
<< pdcontact >>
rect 4 -2 8 6
rect 12 -2 16 6
rect 42 -2 46 6
rect 50 -2 54 6
<< polysilicon >>
rect 9 6 11 9
rect 47 6 49 9
rect 9 -17 11 -2
rect 47 -17 49 -2
rect 9 -24 11 -21
rect 47 -24 49 -21
<< polycontact >>
rect 5 -14 9 -10
rect 43 -14 47 -10
<< metal1 >>
rect -2 11 23 15
rect 36 11 61 15
rect 4 6 8 11
rect 42 6 46 11
rect 12 -10 16 -2
rect 50 -10 54 -2
rect -8 -14 5 -10
rect 12 -14 43 -10
rect 50 -14 70 -10
rect 12 -17 16 -14
rect 50 -17 54 -14
rect 4 -25 8 -21
rect 42 -25 46 -21
rect -2 -29 24 -25
rect 36 -29 62 -25
<< labels >>
rlabel metal1 -2 -29 24 -25 1 GND
rlabel metal1 2 14 19 15 5 VDD
rlabel metal1 21 -14 31 -11 1 OUTPUT
rlabel metal1 -7 -14 -2 -10 3 INPUT
rlabel metal1 36 -29 62 -25 1 GND
rlabel metal1 40 14 57 15 5 VDD
rlabel metal1 59 -14 69 -11 1 OUTPUT
rlabel metal1 31 -14 36 -10 3 INPUT
<< end >>
