magic
tech scmos
timestamp 1725621116
<< error_s >>
rect 5 71 9 72
rect 13 71 17 72
rect 10 65 12 66
rect 5 48 6 63
rect 16 48 17 63
rect 5 45 17 48
rect 13 44 17 45
rect 17 40 18 44
rect 13 35 17 36
rect 17 31 18 35
rect 13 27 17 28
rect 17 23 18 27
rect 10 13 12 14
<< nwell >>
rect 0 42 22 74
<< ntransistor >>
rect 10 16 12 22
<< ptransistor >>
rect 10 45 12 63
<< ndiffusion >>
rect 9 16 10 22
rect 12 16 13 22
<< pdiffusion >>
rect 9 45 10 63
rect 12 45 13 63
<< ndcontact >>
rect 5 16 9 22
rect 13 16 17 22
<< pdcontact >>
rect 5 45 9 63
rect 13 45 17 63
<< psubstratepcontact >>
rect 5 7 9 11
rect 13 7 17 11
<< nsubstratencontact >>
rect 5 68 9 72
rect 13 68 17 72
<< polysilicon >>
rect 10 63 12 65
rect 10 22 12 45
rect 10 14 12 16
<< polycontact >>
rect 6 31 10 35
<< metal1 >>
rect 0 72 22 74
rect 0 68 5 72
rect 9 68 13 72
rect 17 68 22 72
rect 0 66 22 68
rect 5 63 9 66
rect 13 44 17 45
rect 0 31 6 35
rect 17 31 22 35
rect 13 22 17 23
rect 5 13 9 16
rect 0 11 22 13
rect 0 7 5 11
rect 9 7 13 11
rect 17 7 22 11
rect 0 5 22 7
<< m2contact >>
rect 13 40 17 44
rect 13 31 17 35
rect 13 23 17 27
<< metal2 >>
rect 13 35 17 40
rect 13 27 17 31
use my_inverter  my_inverter_0
timestamp 1725621116
transform 1 0 43 0 1 72
box -8 -29 70 15
<< labels >>
rlabel metal1 3 33 3 33 1 in
rlabel metal1 19 33 19 33 1 out
rlabel metal1 11 70 11 70 1 Vdd
rlabel metal1 11 9 11 9 1 GND
<< end >>
